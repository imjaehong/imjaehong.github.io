`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);

    logic [31:0] rom[0:61];

    initial begin
        //rom[x]=32'b func7 _ rs2 _ rs1 _f3 _ rd  _  op
        rom[0] = 32'b0000000_00010_00001_000_00011_0110011;  // add  x3, x1, x2
        rom[1] = 32'b0100000_00010_00001_000_00011_0110011;  // sub  x3, x1, x2
        rom[2] = 32'b0000000_00010_00001_001_00011_0110011;  // sll  x3, x1, x2
        rom[3] = 32'b0000000_00010_00001_101_00011_0110011;  // srl  x3, x1, x2
        rom[4] = 32'b0100000_00010_00001_101_00011_0110011;  // sra  x3, x1, x2
        rom[5] = 32'b0000000_00010_00001_010_00011_0110011;  // slt  x3, x1, x2
        rom[6] = 32'b0000000_00010_00001_011_00011_0110011;  // sltu x3, x1, x2
        rom[7] = 32'b0000000_00010_00001_100_00011_0110011;  // xor  x3, x1, x2
        rom[8] = 32'b0000000_00010_00001_110_00011_0110011;  // or   x3, x1, x2
        rom[9] = 32'b0000000_00010_00001_111_00011_0110011;  // and  x3, x1, x2
    end


    // 하위 2bit 를 없애면 4(2^2)의 배수로 표현이 됨, 4byte 단위로 이동 가능
    assign data = rom[addr[31:2]];

endmodule
